
module bsg_bladerunner_configuration #(parameter width_p=-1, addr_width_p=-1)
(input  [addr_width_p-1:0] addr_i
,output logic [width_p-1:0]      data_o
);
always_comb case(addr_i)
         0: data_o = width_p ' (32'b00000000000000110000011000000010); // 0x00030602
         1: data_o = width_p ' (32'b00000101000000010010000000100000); // 0x05012020
         2: data_o = width_p ' (32'b00000000000000000000000000011100); // 0x0000001C
         3: data_o = width_p ' (32'b00000000000000000000000000100000); // 0x00000020
         4: data_o = width_p ' (32'b00000000000000000000000000001001); // 0x00000009
         5: data_o = width_p ' (32'b00000000000000000000000000001111); // 0x0000000F
         6: data_o = width_p ' (32'b00000000000000000000000000000000); // 0x00000000
         7: data_o = width_p ' (32'b00000000000000000000000000000000); // 0x00000000
         8: data_o = width_p ' (32'b00000000000000000000000000000000); // 0x00000000
         9: data_o = width_p ' (32'b00000111111011001001110100111110); // 0x07EC9D3E
        10: data_o = width_p ' (32'b00000010110001111100010100111100); // 0x02C7C53C
        11: data_o = width_p ' (32'b00000101101100000101011001110100); // 0x05B05674
        12: data_o = width_p ' (32'b00000000000000000000000000000010); // 0x00000002
        13: data_o = width_p ' (32'b00000000000000000000001000000000); // 0x00000200
        14: data_o = width_p ' (32'b00000000000000000000000000001000); // 0x00000008
        15: data_o = width_p ' (32'b00000000000000000000000000001000); // 0x00000008
        16: data_o = width_p ' (32'b00000000000000000000000000100000); // 0x00000020
        17: data_o = width_p ' (32'b00000000000000000000000000100000); // 0x00000020
        18: data_o = width_p ' (32'b00000000000000000000000100000000); // 0x00000100
        19: data_o = width_p ' (32'b00000000000000000000000011001000); // 0x000000C8
   default: data_o = 'X;
endcase
endmodule