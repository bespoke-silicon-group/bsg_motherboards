`ifndef BSG_BLADERUNNER_ROM_PKG
`define BSG_BLADERUNNER_ROM_PKG

package bsg_bladerunner_rom_pkg;

parameter rom_width_gp = 32;
parameter rom_els_gp = 20;

endpackage

`endif
